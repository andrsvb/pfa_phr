----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12.05.2020 13:04:30
-- Design Name: 
-- Module Name: decoder_puntuacion - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

--Traduce las posiciones abstraidas a enteros al array de bits que permite su representación en el display de 7 segmentos.

entity decoder_posicion is
 Port ( 
  posicion_d : in integer range 0 to 2;
  leds : out std_logic_vector (7 downto 0)
  );
end decoder_posicion;

architecture Behavioral of decoder_posicion is

begin

leds <= "11101111" when posicion_d=0 else
        "11111101" when posicion_d=1 else
        "01111111" when posicion_d=2;

end Behavioral;
