----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12.05.2020 13:04:30
-- Design Name: 
-- Module Name: decoder_puntuacion - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

--Aumenta en uno el entero recibido dentro del rango aceptado dando la vuelta si llega el más elevado, 
--este componente se usa para actualizar la posición del personaje del jugador abastraida a un entero.

entity up_pos is
 Port ( 
  posicion_u : in integer range 0 to 2;
  u_posicion : out integer range 0 to 2 
  );
end up_pos;

architecture Behavioral of up_pos is

begin

u_posicion <= 1 when posicion_u=0 else
              2 when posicion_u=1 else
              0 when posicion_u=2;

end Behavioral;
